.TITLE exemplo 01

* ****************************************************************************
*        1   2   3
*        +-@-+-@-+-
*        |   |   |
*        @   @   =
*        |   |
*       (~)  =
*        |
*        =

* ****************************************************************************
*            3   0
*        +-@-+-@-+-
*     2  |   |   |
*        @   @   = 0
*     1  |   |
*       (~)  = 0
*        |
*     0  =

V1    1 0   10V
xdiv1 2 3 0 vdivide
R1    3 0   5K

* The following are the subcircuit definition cards:
*
.subckt vdivide 1 2 3
r1 1 2 10K
r2 2 3 5K
.ends

.op

.end

